library verilog;
use verilog.vl_types.all;
entity tb_arithmetic_unit is
end tb_arithmetic_unit;
